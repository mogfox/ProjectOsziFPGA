-- intADC_tb.vhd

-- Generated using ACDS version 20.1 711

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity intADC_tb is
end entity intADC_tb;

architecture rtl of intADC_tb is
	component intADC is
		port (
			adc_pll_clock_clk      : in  std_logic                     := 'X';             -- clk
			adc_pll_locked_export  : in  std_logic                     := 'X';             -- export
			clock_clk              : in  std_logic                     := 'X';             -- clk
			command_valid          : in  std_logic                     := 'X';             -- valid
			command_channel        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- channel
			command_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			command_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			command_ready          : out std_logic;                                        -- ready
			reset_sink_reset_n     : in  std_logic                     := 'X';             -- reset_n
			response_valid         : out std_logic;                                        -- valid
			response_channel       : out std_logic_vector(4 downto 0);                     -- channel
			response_data          : out std_logic_vector(11 downto 0);                    -- data
			response_startofpacket : out std_logic;                                        -- startofpacket
			response_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component intADC;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal intadc_inst_adc_pll_clock_bfm_clk_clk  : std_logic; -- intADC_inst_adc_pll_clock_bfm:clk -> intADC_inst:adc_pll_clock_clk
	signal intadc_inst_clock_bfm_clk_clk          : std_logic; -- intADC_inst_clock_bfm:clk -> [intADC_inst:clock_clk, intADC_inst_reset_sink_bfm:clk]
	signal intadc_inst_reset_sink_bfm_reset_reset : std_logic; -- intADC_inst_reset_sink_bfm:reset -> intADC_inst:reset_sink_reset_n

begin

	intadc_inst : component intADC
		port map (
			adc_pll_clock_clk      => intadc_inst_adc_pll_clock_bfm_clk_clk,  --  adc_pll_clock.clk
			adc_pll_locked_export  => open,                                   -- adc_pll_locked.export
			clock_clk              => intadc_inst_clock_bfm_clk_clk,          --          clock.clk
			command_valid          => open,                                   --        command.valid
			command_channel        => open,                                   --               .channel
			command_startofpacket  => open,                                   --               .startofpacket
			command_endofpacket    => open,                                   --               .endofpacket
			command_ready          => open,                                   --               .ready
			reset_sink_reset_n     => intadc_inst_reset_sink_bfm_reset_reset, --     reset_sink.reset_n
			response_valid         => open,                                   --       response.valid
			response_channel       => open,                                   --               .channel
			response_data          => open,                                   --               .data
			response_startofpacket => open,                                   --               .startofpacket
			response_endofpacket   => open                                    --               .endofpacket
		);

	intadc_inst_adc_pll_clock_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => intadc_inst_adc_pll_clock_bfm_clk_clk  -- clk.clk
		);

	intadc_inst_clock_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => intadc_inst_clock_bfm_clk_clk  -- clk.clk
		);

	intadc_inst_reset_sink_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => intadc_inst_reset_sink_bfm_reset_reset, -- reset.reset_n
			clk   => intadc_inst_clock_bfm_clk_clk           --   clk.clk
		);

end architecture rtl; -- of intADC_tb
