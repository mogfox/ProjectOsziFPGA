------------------------------------------------------------------------------------
--Project : DIC 3BHEL 
--Author  : Gr�bner
--Date    : 15/05/2018
--File    : DE10_Lite_const_pkg.vhd
--Design  : Terasic DE10 Board
------------------------------------------------------------------------------------
-- Description: Single Pulse Generation for Pushbutton
------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;

--=======================================================================================================
entity pulse_gen is
  port (
        RESET_n   :  in std_logic;
        CLK_50MHz :  in std_logic;
        BUTTON_in :  in std_logic;
        PULSE_out : out std_logic
       );
end pulse_gen;
--=======================================================================================================

--&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
architecture rtl of pulse_gen is
  --=====================================================================================================
  type state_type is (ST_IDLE, ST_PULSE, ST_WAIT); 
  signal state : state_type;
  --=====================================================================================================
begin
  --=====================================================================================================
  PulseGen: process(CLK_50MHz, RESET_n)
  begin
    if (RESET_n = '0') then
      state     <= ST_IDLE;
      PULSE_out <= '0';
    elsif (CLK_50MHz'event and CLK_50MHz = '1') then
      case state is
        -------------------------------------------------------------------------------------------------
        when ST_IDLE  =>
          if (BUTTON_in = '1') then
            state     <= ST_PULSE;
            PULSE_out <= '1';
          end if;
        -------------------------------------------------------------------------------------------------
        when ST_PULSE =>
          PULSE_out <= '0';
          if (BUTTON_in = '1') then
            state <= ST_WAIT;
          else
            state <= ST_IDLE;
          end if;
        -------------------------------------------------------------------------------------------------
        when ST_WAIT  =>
          if (BUTTON_in = '0') then
            state <= ST_IDLE;
          end if;
        -------------------------------------------------------------------------------------------------
        when others => NULL;
        -------------------------------------------------------------------------------------------------
      end case;
    end if;
  end process PulseGen;
  --=====================================================================================================
end rtl;
--&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
